LIBRARY ieee;

USE ieee.std_logic_1164.ALL;


ENTITY ALU IS
PORT
(
	input1: IN std_logic_vector(15 DOWNTO 0);
	input2: IN std_logic_vector(15 DOWNTO 0);
	output: OUT std_logic_vector(15 DOWNTO 0)
);
END ALU;

ARCHITECTURE Struct OF ALU IS
BEGIN
END Struct;